module moduleName (
    ports
);
    // TODO
endmodule