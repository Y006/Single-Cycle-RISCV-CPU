module tb_memory;

memory U_memory
(

);

initial begin

end

endmodule