module memory (
    input  [0 :4] I_address,
    input         I_mem_wirte_en,
    input  [31:0] I_data,
    output [31:0] O_data
);


endmodule